module test04(
    input  clk,
    output dout
);

endmodule
