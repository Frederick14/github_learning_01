module test04(
    input clk
);

endmodule