module test04(

);

endmodule